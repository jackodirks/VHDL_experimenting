library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library vunit_lib;
context vunit_lib.vunit_context;
context vunit_lib.vc_context;

library src;
use src.mips32_pkg;

entity mips32_coprocessor_zero_tb is
    generic (
        runner_cfg : string);
end entity;

architecture tb of mips32_coprocessor_zero_tb is
    constant clk_period : time := 20 ns;

    signal clk : std_logic := '0';
    signal rst : std_logic := '0';

    signal address_from_controller : natural range 0 to 31 := 0;
    signal address_from_pipeline : natural range 0 to 31 := 0;

    signal write_from_controller : boolean := false;
    signal write_from_pipeline : boolean := false;

    signal data_from_controller : mips32_pkg.mips32_data_type := (others => '0');
    signal data_from_pipeline : mips32_pkg.mips32_data_type := (others => '0');

    signal data_to_controller : mips32_pkg.mips32_data_type;
    signal data_to_pipeline : mips32_pkg.mips32_data_type;

    signal cpu_reset : boolean;
    signal cpu_stall : boolean;

begin

    clk <= not clk after (clk_period/2);

    main : process
    begin
        test_runner_setup(runner, runner_cfg);
        while test_suite loop
            if run("cpu reset is true before first rising edge") then
                wait until rising_edge(clk);
                check(cpu_reset);
            elsif run("data_to_controller address 0 reads as 1 before first rising edge") then
                address_from_controller <= 0;
                wait until rising_edge(clk);
                check(X"00000001" = data_to_controller);
            elsif run("data_to_controller address 5 reads as 0 before first rising edge") then
                address_from_controller <= 5;
                wait until rising_edge(clk);
                check(X"00000000" = data_to_controller);
            elsif run("data_to_pipeline address 0 reads as 1 before first rising edge") then
                address_from_pipeline <= 0;
                wait until rising_edge(clk);
                check(X"00000001" = data_to_pipeline);
            elsif run("data_to_pipeline address 5 reads as 0 before first rising edge") then
                address_from_pipeline <= 5;
                wait until rising_edge(clk);
                check(X"00000000" = data_to_pipeline);
            elsif run("Writing 0 to address 0 from data_from_controller drops cpu_reset") then
                wait until falling_edge(clk);
                address_from_controller <= 0;
                data_from_controller <= (others => '0');
                write_from_controller <= true;
                wait until falling_edge(clk);
                check(not cpu_reset);
            elsif run("Read after write from controller returns last written data") then
                wait until falling_edge(clk);
                address_from_controller <= 0;
                data_from_controller <= (others => '0');
                write_from_controller <= true;
                wait until falling_edge(clk);
                write_from_controller <= false;
                wait until rising_edge(clk);
                check(X"00000000" = data_to_controller);
            elsif run("Writing 0 to address 5 from data_from_controller keep cpu_reset high") then
                wait until falling_edge(clk);
                address_from_controller <= 5;
                data_from_controller <= (others => '0');
                write_from_controller <= true;
                wait until falling_edge(clk);
                check(cpu_reset);
            elsif run("Read from pipeline after controller write returns last written data") then
                wait until falling_edge(clk);
                address_from_controller <= 0;
                data_from_controller <= (others => '0');
                write_from_controller <= true;
                address_from_pipeline <= 0;
                write_from_pipeline <= false;
                wait until falling_edge(clk);
                write_from_controller <= false;
                wait until rising_edge(clk);
                check(X"00000000" = data_to_pipeline);
            elsif run("Writing 0 to address 0 from data_from_pipeline drops cpu_reset") then
                wait until falling_edge(clk);
                address_from_pipeline <= 0;
                data_from_pipeline <= (others => '0');
                write_from_pipeline <= true;
                wait until falling_edge(clk);
                check(not cpu_reset);
            elsif run("Writing 0 to address 5 from data_from_pipeline keeps cpu_reset high") then
                wait until falling_edge(clk);
                address_from_pipeline <= 5;
                data_from_pipeline <= (others => '0');
                write_from_pipeline <= true;
                wait until falling_edge(clk);
                check(cpu_reset);
            elsif run("Writing 2 to address 0 disables reset, enables stall") then
                wait until falling_edge(clk);
                address_from_controller <= 0;
                data_from_controller <= X"00000002";
                write_from_controller <= true;
                wait until falling_edge(clk);
                check(not cpu_reset);
                check(cpu_stall);
            elsif run("Only bits 0 and 1 are writable") then
                wait until falling_edge(clk);
                address_from_pipeline <= 0;
                data_from_pipeline <= (others => '1');
                write_from_pipeline <= true;
                wait until falling_edge(clk);
                write_from_pipeline <= false;
                wait until rising_edge(clk);
                check(data_to_pipeline = X"00000003");
            elsif run("rst resets") then
                wait until falling_edge(clk);
                address_from_controller <= 0;
                data_from_controller <= X"00000002";
                write_from_controller <= true;
                wait until falling_edge(clk);
                write_from_controller <= false;
                rst <= '1';
                wait until falling_edge(clk);
                check(cpu_reset);
                check(not cpu_stall);
            end if;
        end loop;
        wait until rising_edge(clk);
        wait until falling_edge(clk);
        test_runner_cleanup(runner);
        wait;
    end process;

    test_runner_watchdog(runner,  1 us);

    coprocessor_zero : entity src.mips32_coprocessor_zero
    port map (
        clk,
        rst,
        address_from_controller,
        address_from_pipeline,
        write_from_controller,
        write_from_pipeline,
        data_from_controller,
        data_from_pipeline,
        data_to_controller,
        data_to_pipeline,
        cpu_reset,
        cpu_stall
    );
end architecture;
